LIBRARY  IEEE;                                              
USE IEEE.STD_LOGIC_1164.ALL;				
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
ENTITY  mq_clock_top IS
PORT (CLKK: IN  STD_LOGIC;
	  RST1: IN  STD_LOGIC;
	  SET_H: IN  STD_LOGIC;
	  SET_M: IN  STD_LOGIC;
	  LED2H,LED1H,LED2M,LED1M,LED2S,LED1S,led2z,led2c: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
	  --LED2S HEX1 秒（十位）     LED1S HEX0 秒（个位）
	  --LED2H HEX5 小时（十位）    LED1H  HEX4 小时（个位）
     --LED2M HEX3 分钟（十位）	  LED1M  HEX2 分钟（个位）
	  LIGHT_O: OUT  STD_LOGIC_VECTOR(7 DOWNTO 0));
END  ENTITY  mq_clock_top;		
ARCHITECTURE  FOUR  OF  mq_clock_top IS
COMPONENT  FENPIN                         
PORT (CLK50: IN  STD_LOGIC;
	 				CLK1HZ: OUT  STD_LOGIC;
	 				CLKZOU: OUT  STD_LOGIC_VECTOR(1 DOWNTO 0));
END  COMPONENT;
COMPONENT  SETTIME
PORT (CLK: IN  STD_LOGIC;RST: IN  STD_LOGIC;
	  				SETH: IN  STD_LOGIC;SETM: IN  STD_LOGIC;
	HOUR2,HOUR1,MIN2,MIN1,SEC2,SEC1: BUFFER  STD_LOGIC_VECTOR(3 DOWNTO 0);
	             ZOUMA: OUT  STD_LOGIC);
END  COMPONENT;
COMPONENT  LED
PORT (H2,H1,M2,M1,S2,S1: IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
	 LEDH2,LEDH1,LEDM2,LEDM1,LEDS2,LEDS1:  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0));
END  COMPONENT;
COMPONENT  ZOUMADENG
PORT(ZOU_MA: IN  STD_LOGIC;
	          CLKZ: IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
	          LIGHT: OUT  STD_LOGIC_VECTOR(7 DOWNTO 0));
END  COMPONENT;
SIGNAL  a,ss: STD_LOGIC;
SIGNAL  b,c,d,e,f,g :STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL  tt: STD_LOGIC_VECTOR(1 DOWNTO 0);
BEGIN
led2z<="1111111";
led2c<="1111111";													
U1: FENPIN PORT MAP(CLK50=>CLKK,CLK1HZ=>a,CLKZOU=>tt);
U2:SETTIME PORT MAP(CLK=>a,RST=>RST1,SETH=>SET_H,SETM=>SET_M,HOUR2=>b,HOUR1=>c,MIN2=>d,MIN1=>e,SEC2=>f,SEC1=>g,ZOUMA=>ss);
U3: LED PORT  MAP(H2=>b,H1=>c,M2=>d,M1=>e,S2=>f,S1=>g,LEDH2=>LED2H,LEDH1=>LED1H,LEDM2=>LED2M,LEDM1=>LED1M,LEDS2=>LED2S,LEDS1=>LED1S);
U4: ZOUMADENG  PORT MAP(CLKZ=>tt,ZOU_MA=>ss,LIGHT=>LIGHT_O);
END  ARCHITECTURE  FOUR;
