LIBRARY  IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY  ZOUMADENG  IS
PORT(ZOU_MA: IN  STD_LOGIC;
	 CLKZ: IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
	 LIGHT: OUT  STD_LOGIC_VECTOR(7 DOWNTO 0));
END  ENTITY  ZOUMADENG;
ARCHITECTURE  one  OF  ZOUMADENG  IS
BEGIN
PROCESS(ZOU_MA,CLKZ)  BEGIN
IF  ZOU_MA='1'  THEN 							
		          CASE  CLKZ  IS
		             WHEN "00"=>LIGHT<="01010101";			
		             WHEN "01"=>LIGHT<="10101010";
		             WHEN "10"=>LIGHT<="00000000";
		             WHEN "11"=>LIGHT<="11111111";
		          END  CASE;
ELSIF  ZOU_MA='0'  THEN
	            LIGHT<="00000000";
END  IF;
END  PROCESS;
END  one;