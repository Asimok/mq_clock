LIBRARY  IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
ENTITY  LED  IS

PORT (H2,H1,M2,M1,S2,S1: IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
LEDH2,LEDH1,LEDM2,LEDM1,LEDS2,LEDS1:OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END  ENTITY LED;
ARCHITECTURE  one  OF  LED  IS
BEGIN
PROCESS(H2)  BEGIN									
	    CASE  H2  IS
		       WHEN "0000"=>LEDH2<="1000000"; 
		       WHEN "0001"=>LEDH2<="1111001"; 
		       WHEN "0010"=>LEDH2<="0100100"; 
		       WHEN  OTHERS=>NULL;
	    END  CASE;
END  PROCESS;
PROCESS(H1)  BEGIN								  
	    CASE  H1  IS 
		       WHEN "0000"=>LEDH1<="1000000"; 
		       WHEN "0001"=>LEDH1<="1111001"; 
		       WHEN "0010"=>LEDH1<="0100100"; 
		       WHEN "0011"=>LEDH1<="0110000"; 
		       WHEN "0100"=>LEDH1<="0011001"; 
		       WHEN "0101"=>LEDH1<="0010010"; 
		       WHEN "0110"=>LEDH1<="0000010";
		       WHEN "0111"=>LEDH1<="1111000"; 
		       WHEN "1000"=>LEDH1<="0000000"; 
		       WHEN "1001"=>LEDH1<="0010000";
		       WHEN  OTHERS=>NULL;
	   END  CASE;
END  PROCESS;
PROCESS(M2)  BEGIN									
	   CASE  M2  IS 
		      WHEN "0000"=>LEDM2<="1000000"; 
		      WHEN "0001"=>LEDM2<="1111001"; 
		      WHEN "0010"=>LEDM2<="0100100"; 
		      WHEN "0011"=>LEDM2<="0110000"; 
		      WHEN "0100"=>LEDM2<="0011001"; 
		      WHEN "0101"=>LEDM2<="0010010"; 
		      WHEN  OTHERS=>NULL;
	    END  CASE;
END  PROCESS;
PROCESS(M1)  BEGIN								   
	        CASE  M1  IS 
		       WHEN "0000"=>LEDM1<="1000000"; 
		       WHEN "0001"=>LEDM1<="1111001"; 
		       WHEN "0010"=>LEDM1<="0100100"; 
		       WHEN "0011"=>LEDM1<="0110000"; 
		       WHEN "0100"=>LEDM1<="0011001"; 
		       WHEN "0101"=>LEDM1<="0010010"; 
		       WHEN "0110"=>LEDM1<="0000010";
		       WHEN "0111"=>LEDM1<="1111000"; 
		       WHEN "1000"=>LEDM1<="0000000"; 
		       WHEN "1001"=>LEDM1<="0010000";
		       WHEN  OTHERS=>NULL;
	        END  CASE;
END  PROCESS;
PROCESS(S2)  BEGIN									 
	       CASE  S2  IS 
		      WHEN "0000"=>LEDS2<="1000000"; 
		      WHEN "0001"=>LEDS2<="1111001"; 
		      WHEN "0010"=>LEDS2<="0100100"; 
		      WHEN "0011"=>LEDS2<="0110000"; 
		      WHEN "0100"=>LEDS2<="0011001"; 
		      WHEN "0101"=>LEDS2<="0010010"; 
		      WHEN  OTHERS=>NULL;
	       END  CASE;
END  PROCESS;
PROCESS(S1)  BEGIN								
	       CASE  S1  IS 
		      WHEN "0000"=>LEDS1<="1000000"; 
		      WHEN "0001"=>LEDS1<="1111001"; 
		      WHEN "0010"=>LEDS1<="0100100"; 
		      WHEN "0011"=>LEDS1<="0110000"; 
		      WHEN "0100"=>LEDS1<="0011001"; 
		      WHEN "0101"=>LEDS1<="0010010"; 
		      WHEN "0110"=>LEDS1<="0000010";
		      WHEN "0111"=>LEDS1<="1111000"; 
		      WHEN "1000"=>LEDS1<="0000000"; 
		      WHEN "1001"=>LEDS1<="0010000";
		      WHEN  OTHERS=>NULL;
	     END  CASE;
END  PROCESS;
END  ARCHITECTURE  one;